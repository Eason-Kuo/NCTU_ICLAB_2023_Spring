`ifdef RTL
`define CYCLE_TIME 5
	`define RTL_GATE
`elsif GATE
`define CYCLE_TIME 5
	`define RTL_GATE
`elsif CHIP
`define CYCLE_TIME 5
    `define CHIP_POST 
`elsif POST
`define CYCLE_TIME 5
    `define CHIP_POST 
`endif

`define CYCLE_TIME_DATA 31.7

`ifdef FUNC
`define PAT_NUM 836
`define MAX_WAIT_READY_CYCLE 2000
`endif
`ifdef PERF
`define PAT_NUM 836
`define MAX_WAIT_READY_CYCLE 100000
`endif


`include "../00_TESTBED/MEM_MAP_define.v"
`include "../00_TESTBED/pseudo_DRAM_data.v"
`include "../00_TESTBED/pseudo_DRAM_inst.v"

module PATTERN(
    			clk,
			  rst_n,
		   IO_stall,


         awid_s_inf,
       awaddr_s_inf,
       awsize_s_inf,
      awburst_s_inf,
        awlen_s_inf,
      awvalid_s_inf,
      awready_s_inf,
                    
        wdata_s_inf,
        wlast_s_inf,
       wvalid_s_inf,
       wready_s_inf,
                    
          bid_s_inf,
        bresp_s_inf,
       bvalid_s_inf,
       bready_s_inf,
                    
         arid_s_inf,
       araddr_s_inf,
        arlen_s_inf,
       arsize_s_inf,
      arburst_s_inf,
      arvalid_s_inf,
                    
      arready_s_inf, 
          rid_s_inf,
        rdata_s_inf,
        rresp_s_inf,
        rlast_s_inf,
       rvalid_s_inf,
       rready_s_inf 
    );

//---------------------------------------------------------------------
//   PORT DECLARATION          
//---------------------------------------------------------------------
parameter ID_WIDTH=4, DATA_WIDTH=32, ADDR_WIDTH=32, DRAM_NUMBER=2, WRIT_NUMBER=1;

output reg			  clk,rst_n;
input				IO_stall;

// axi write address channel 
input wire [WRIT_NUMBER * ID_WIDTH-1:0]        awid_s_inf;
input wire [WRIT_NUMBER * ADDR_WIDTH-1:0]    awaddr_s_inf;
input wire [WRIT_NUMBER * 3 -1:0]            awsize_s_inf;
input wire [WRIT_NUMBER * 2 -1:0]           awburst_s_inf;
input wire [WRIT_NUMBER * 7 -1:0]             awlen_s_inf;
input wire [WRIT_NUMBER-1:0]                awvalid_s_inf;
output wire [WRIT_NUMBER-1:0]               awready_s_inf;
// axi write data channel 
input wire [WRIT_NUMBER * DATA_WIDTH-1:0]     wdata_s_inf;
input wire [WRIT_NUMBER-1:0]                  wlast_s_inf;
input wire [WRIT_NUMBER-1:0]                 wvalid_s_inf;
output wire [WRIT_NUMBER-1:0]                wready_s_inf;
// axi write response channel
output wire [WRIT_NUMBER * ID_WIDTH-1:0]         bid_s_inf;
output wire [WRIT_NUMBER * 2 -1:0]             bresp_s_inf;
output wire [WRIT_NUMBER-1:0]             	  bvalid_s_inf;
input wire [WRIT_NUMBER-1:0]                  bready_s_inf;
// -----------------------------
// axi read address channel 
input wire [DRAM_NUMBER * ID_WIDTH-1:0]       arid_s_inf;
input wire [DRAM_NUMBER * ADDR_WIDTH-1:0]   araddr_s_inf;
input wire [DRAM_NUMBER * 7 -1:0]            arlen_s_inf;
input wire [DRAM_NUMBER * 3 -1:0]           arsize_s_inf;
input wire [DRAM_NUMBER * 2 -1:0]          arburst_s_inf;
input wire [DRAM_NUMBER-1:0]               arvalid_s_inf;
output wire [DRAM_NUMBER-1:0]              arready_s_inf;
// -----------------------------
// axi read data channel 
output wire [DRAM_NUMBER * ID_WIDTH-1:0]         rid_s_inf;
output wire [DRAM_NUMBER * DATA_WIDTH-1:0]     rdata_s_inf;
output wire [DRAM_NUMBER * 2 -1:0]             rresp_s_inf;
output wire [DRAM_NUMBER-1:0]                  rlast_s_inf;
output wire [DRAM_NUMBER-1:0]                 rvalid_s_inf;
input wire [DRAM_NUMBER-1:0]                  rready_s_inf;
// -----------------------------





//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
Ff4XRvHaSSXYDl1lyydTyCM/GlEEh1kJmDTYFyT4ceZCyL+W6HwB1pjzqx8cU/L3
o5uKBIorw3ZzJjgjJL3jZ/MOgnIOoJnZt8YnxgIUfh7XSHnQ2B7PJs9eX2dizD5H
Vo8gnkmnGKxj2aMO2bLBUDqFblMVij7pwHNmwh3+UQBw2H9tU2innD5VOmjxq8Ow
9JoPp6zvXjdhgMN+X+ad4I653b542vVUbSYwBRh+z7h7N1vSzkH98LWfb6BDF+4D
WirsbmE09khgN8cMj3UVc+EL2L3bzeN7Wr8vZJISfxN37jaLyBJkugq2yb5p0o7U
9Rh9wvHA4enRHVfpotZ7CQ==
//pragma protect end_key_block
//pragma protect digest_block
xr64PRJr7p/kx/SRzvrONcgj5Sc=
//pragma protect end_digest_block
//pragma protect data_block
KYVc747GPqatTGzqDWB3pmg0JG4xBqu9gwcHzlZ1VFl1oFrDhn6eoWpdibgNIyse
4WapMWUANoTiQj+6mqyitWT3JvTCuQK8ffj2doTTqaG9tdqOM2pbf08JHRfiTWMj
t56svmGFFofEmnDVfctKURRH91+6B++DuQ69Cb7I/Naq53nGEOkPYTxUEVmaaxuI
8Qt+jOANijBFL7LEN8gSMwK8UsApY9uSakiknZOoUCiEetp0lGjIwzWtVyRT085y
mQ696bOrjjopTF/h12yIBaGigDqBf42Yq4HB8rwkW9uKyur9uPJ5YTR5bUJemE90
3kexbIcyNanLmm1aNaoMx/lmVrZ0rUPBkhuJzNV/0e6GXGGFJzpeR6uMDoTfGOl3
WaAibfxKfq9/qNxYcwi3ifM6u6HEi47OAbrpDD/nOA+sSk4Uhyvq8K2mvyDAigso
iOGCRtK/BmlSlI/r0iGCXiTXpmCzihr5lJ60t5h5XcVYA+YhkhyrlD8t0UlkqfbK
oS3/YlNRNgsFQf8qj1QViJ3n2gT5cskZsfumFUPJcvfut+c3NQzXkxAV3woT6tSg
CRi3aFNblyGvW+noZ6ZYOttHBN2/cX2MbIwEJRpZIN96GhICGig0rILWwCAuN+BG
v0tr6VLv5JsVrrfI5EtGF8R/KJmZXLTifjZG3+IfxyKAA2S+HMz+lTuXFvaO0lRZ
COnpMYqkF4WyxQaF9uKMuXHMqoLB2cFdi2AoJFeNxdmnRQiNYzzZsMv27i1hJZtP
o/DPVevm6BmH7xSpW88wxWo9f12uwXHyZc+BiozB2eiNnSVeMtZFcPqONoeu36ZL
Nyh2jS2LqMYsAIpvj2BTmu8fsRUTHJcCH1KuscFZ+dm51P1a5gvbWRlvAScy6BYi
BfDxPUiVrizS1M2SvLF3DTSz4Bf9EEircXyMCaLOz+DNx/S3htXIKR6UbmPx4AmR
7Vp0/bw77O70nD+Cxum7ZJ2z3MwbRFj7M9Ny1m/88MJ+NdvtVZ9JD+n9Z3eVk7RS
kKQUiNNRPRTDgvNvTgSV8qJ5ql2YyljwCHasJRUUQzjKu5/dz/kz95UufdD0dsOR
lIK5xfSssKpNBD5ijdlZddBPpVcTijLvC06DH3x7dQIjVp0N8tDZneNGHWhL/9eX
gvmOjihgVjIp7E4JKodwhUmlfNsnByPYOvQvxPcdgiQwvpC7xZBdVHHasAcz/OmS
L1TJjUc4O+6NbGsgm90kdlv7M9S9P08Wqz3opZQ2lahB21RIVeIvYJRUALpdc0Z8
WK5JDj9eZNy5Cphpw7CEfntClWSfGufnH7u/7ZNdudkRMOOgqzmu5jbJhtItttmd
okkd/dpstWJau6DuPxYivy4Hi6H796i/1JkXKHTf1wB4vVpFfPnL9qBc1NQ34gP7
x4zvvxKOhxRpEeMz3+ZmlYByPzMdXGEknslPLCU0FHbGLRi/c6MHPRyygzKXpuQO
XVLKgGWTNS9IrrkJzGWiKs5IcynkBkzODPr/E1c8re+kz/HRCROOGlvJOVkkF2Q6
ipG3be4ojFUelKWhcHQZlIVvaKjeshWwTPCunFYLHnUtf4gYDD9lGX6wP1AiZzYM
yOUXM61kXAHn6K6hTQxto6E+SxfXzfPZgRzcADZSJJmUMyz43ikBRlSYhSkcJXzZ
diU/YaXab7NRhGHGQYZlMKtSFWdngHq7t2aKyk2Ezm91emsUlTTGzFRe9BqqvQGA
wqODwNPO04tjWug2vzIT9PzAPOOljGX8HS2s/EM7o2p4vriuaIZCqV0sfnT4sRcb
3yjwCTntRRmoEESAB4zuKYntbE4nHkVUF45NjID93EtHeUi76EZMvVU9lVZKArjf
KUj2Wajaxi0ITS3WoyvTHqcw/TQSJgHYe9U1XIp10K6c6A6760IBuTwhfuA+hChq
PJfJIOkvL4Yz5xlrXWJ74AETKY3iG6l/czn1r9KPC3qOzRECONpPvU8ok5N7oR1w
nPU+5XZzaW/mVpw5UKV/EjJ36ddyd4cQNzdMocO719hpNMLCCOCO+Y5qPLR0Tzs7
/0avpU0xeNDHC+RIYCeelx6vQbcCOYKnIrBXHKktPYytl3zOeKpf+CIBKZtxeTLP
AUO39ugllgVH9OjcG2G7I0y5EwzC/PbV7LiWpdASvQ7UPWf+En3Ttkju82nobqnO
cRuu/D48SZrmXqHVvrtG7+LWi8MRXAJvuiIfcNliy9paRGd1pd2SOmVrl+V9rHMx
+Hswh5ph/7dA5V3eNU4exl2hddOXyy0z/LhKpBvIZfVNWPpafrQ5UiKi2qG6RQtX
9FDrXQJ5Y9y+pAk6WIEuRFJsLHhLAWxxbP1KqPdUF5VabrYnDE81NuXeSSSeRbx1
O1QxQCY91kwhHRXlJzCrqLKgAkXHk+N+zuRfmsHaDivHJirNr8MfNa5jCJYSbZ1K
3+V0UCrdENUNZG3zXwPryRx4FlwWD44aULGG8q0R31V8CEorceYtdMTrbMYlAWDJ
c2uUzwH11aUEILbVsHnCzOnoqQowKxGAWJT0pUKyu5m7yPN23Rq+f8lasyyqVaG9
S+ie4EwFtqWXCL2L2OFqyqeISKsEIE4ER0IZtKj6wnEhy/2oI5nlOPY+vCQfIUa/
iNe34G7s8AoJeYypDiPbzKX15MZ1D9U80dMVE7gT9MClDWoYirB9oJ8EHh/vGDio
0ZBF5PAep0aA0aNbjaV6wJftNJ7LTtDnjMSABN2Aef0UT2KZ7pmG/F6ZPiC+Kqi9
sXqnNMNThZb5orZBAS4qkVMTwGY7GRaNcz/yDCfHhWOwLFeffbHiLWDMLZK41TdC
KnUxNYzHNxbjX17hPEhdiFjqIaHBZjMj5YH0lKkzxTZWIe7XoPtQUe6bUnyoBrkr
Pahx2tn2huFffaMX+2lQsIs6EcETEWhaxaSkIXD1GAdtsfTbEZb2STXlJJNHgnno
wLhoIoiaMKe+PIe2EWHqR0zY+iN8fQH5y9+kHOcHdJIMNqaGdeqM33ON5qFjFGsZ
UGgP23+SeWblR0CsbmDgIlywbDYyS/P0VZ462CaslTjoPSqANdUxaYBaG/0jRGwt
6NcqfBbEvDY1YnZEzhAV27SchjV+KqMk68lxTMmJesFBUgm4KNdWMoQ6r4D6FpbU
0I19+EVF7XGkwwWaRXEZJkcV37hu9NEAOWhdhp67Ox6agmcxRq/axX8/zkz0mRix
SA8Q3AkWfUE/JcBy4HSQsCa2bPEeOJgr7hWUjXCxemCMU6sdwpq0gEGJCxoAA52N
IRrhq+zBQYFO66Hj16odafgjIqab6XyTxkwCLus0AWM7JIiKnKGalZn70v1qTHF/
yPOWbj+XZBTUcPNlJT8ADvZdW7fYB2xQ4VFy/xw31hSl9VYI1WngoZjLcPSjncp2
4Uq0hxta8Rt4mOzADzux4r4k3KEL0e6CtqjiYxYqBK+9XT/WIScjYojQmvXehjtG
Ra6MvPSPfGb9Q2asdfH3kVq9/UFHMT02esLzbSa7iYpAU7HLua3aIR5nRrs8BD5L
rggjCAKgqQL+Oc4I9TTXBiY4ABLj5dOmTw1I0W8eBPDMGY9YTbZVvVgd1aPIrsdU
u46yPmu1uZ2HKVFyuGUeATy4iJS5/mhFhWexhXk3NSPTyClwUuveo93d6gTB3H72
uv7AHahHf6PQA4hreb9H0DWq7AGlxB5cBgTWFfCe8lH7J85NCXT4nCmMgnsCfuMB
8VGlo1KwL066ph8cv7b7SpxQwZ7TvVFFqUybFoxNejnNhsmHxtoHlpJQZ9DF7I1m
FuNjhpkYvfFiyGGYm2vutrVaD96bGoeXoCZGt3IZts1WKkBiD48zjg/YAuBxe5Vq
S2JN5XMe2dpqlCOFSAE9LU3bStQPKvqvJIA6FRx/99s8Rq1B12bhsVlmMzmUyC81
6XzPH6U9CG56CWIoG9/poTOb+eubmlhe12h1MO34hyhJcwRsMF19bQLTCO3u4DUS
7CHr9wuq7q4l0ZJXvkRliK3cyIqDERY+Wz82/iEAoW37wzCaiQtQTnTMRzPaRuYS
j8UIcudtflpff3riHEoQT73AxOmjTIFiqrejP8Ku9YgKvIWKh+hI5e8hVS9lmdlJ
D/Nc4kL8d/380MYEaE0K6I/sxyPAXPaPd1U89N09myp3chEbbp68WkOYpcpChhgl
BSMf1wqueyFFRETc2QsOqFJg8Qemsx5NejfCvQ+w1YBKl9Zfq9BC/eD74Zb1VqQ5
XeyVq64vIREixqKTe2/O1e4C9MvFHprYP9xqPi83DPdJL3yd09MyugJ5pC7IQYMP
suFxOnYTnFHHfkwF3Czl75KnvgqoI0mq8QWTeekBcE3HSwYlTC6JvZ30+qw9pTlv
nSmi+japzu+DVE+lV32H5XT/xprXXLwbuVIhhlZe9/IuIjYzr2ocw1OA6s//BlNz
shzaY9sUQbPlTY/2aMqfNr+FB73pBPVyjewRG/aEWEwPYLQxbHWx3wuFW6CL9F9g
wT8rW4YEmf5S7hux00yIxH59EaaMUKedTGa8CEVYjzDagXyx4cwc/Wv9WAbbYpzJ
i2Cpz5ksYNF8Pzkjrs5c3F+uD389bkQiZ74F9u7wLW0+9OWaPgCnLdHlXUH1SZEz
I+o4LeHkvNl8nc6Xl+A5BBpvOj2wnRaxOwaefO0HB1vQ/4rt3Ssj4g09hhlg2PRn
l6SgqXF6a2gPwUssYPxcoRLYlA/vSjWignytJ2SOUvihwt07YeMDxZ80asz9gu/b
68c/ZLrTSJHqOaSZIw2DvKk7bYSKzZmKXEU1Rq6etYuA1ghQqYLAzIMvGbqIWhkW
AbERycOQDylvk1ohs7Wx40bT4qb26BUfJO6QOceMDNMkxxCZxKgcfikd5ZMbeJNd
8dI1sEMMBvOmC3MumoaVIVZZVh7dPAhhu/OHhjs4NuNEivb8SxTviOJQVcqGUXRa
1gEgr53JbSNm+TEzfhu45HufOKbKQyxwG0HaUelyrT+YjAOopAi+tBkz1IRn32KV
bO2vjT8xfv7QW28qt5na3R4q4v4N1khkGGx+ztvwbqe09lFF50aaHr8PEg4dd+kD
qYXar/OKRSGcTAu7QzwAJlCmtNrizJfhq4R9H1MxIt9r1xg9ttsO09Bg5Ai6m20s
VG24pT6O2lUfiQ1J69ExwNVDXFEkWaynGig36Fj5WR4AQ3RzwzILRQtvWPK+lS9A
gvfA8BWobZhOkeJPMY0lIb+UYEzHL+YZjpgKtjlRGs9QVQEaE44+ohCiZ3kDcLed
2vYj4q036yOGIQz5RT410N0omsWa0vcsNppzKWOF8tpKCBtqQ7QUrLp8bygFHX15
fW0mro7mtVRUrdVQnA7KS27fdndNgfY8cFyxKd79TIIDHXqSaE2sRakPr9dX7ny7
QSPtxVsYjs2Wos7tRtK+MfzhfM08N14Bqb2y8UCdYoflpQceJJzAp1BEnymL+9GQ
+5LXmjxXZy+7NKBj14BsQintAnC4VZrgvy7kUCvbCBawBpeTBYt9pOSFI4H0jPRP
O5OtkLDVj90KU8eDzz3KsGvf9KTHLVKuaTlMUr2VOW9TFghIBdYu34pCsMDQ9xjS
nJr40R9yK8+RYaxJiN/pVRXQm3bH610Moy0rChbsJ06772Qb7wHpBqFPQ+qezEAM
qv6//NJk9KrdtLsDWZp9npnI3+IPRCwASM3ScJ2OvGGnJhtz7HpbAu780MjNUUGN
TjgAjN1O90luyQ9M8VGXwQmjZqlHNNY2kUpfSiFXNThzaP4K8qYjZCpcaRzz+W+X
Iu/leS2wLB8fuOj+1jmmTLu2/FfGOf0AgQGJ6YHQJkAimqd3WkB7DQrXwEA6Dm/g
8mpztfYMVqQU5A1jbzs+UnDIswoF/Bzp3BcBMo/NP1WJxP4UYAFFEVYKKT/EI12P
tAFcf0Yvnjc14p7dG7nPuywMpGtvk8IA4x+2nqSdhm7clalfRK0eZBffeUN7LE9i
otq34wF1YPf731a/iysuzsgh/EeRbPaNNvJ2WanBxt7bqbtVZZB+U9sm9jKEXm/I
vajKRgacS1k3knZpH8fZFtEYoGHGy8QGSNKzl0+4l5O3kgNKqGvxFyf6/Q0NcjBV
gqLG6HTeT8goZMtEDeQkTag6l/T5JbQnUW7gH1iZFkiISAFLTcGg6ll09rvgDRzQ
ex0SfCYviqFYJQe89qwFJgNMzl+LfveE9wbeuTjOH8gafHUt4UMdJRGNFvPEJs2G
YRb1uNo7WXBDTEL20pKflWQmGUtVtHsG23dLmyQPNF7JZvdI61AeJNwApk9UOSNK
2dUrq1TZuKzYxEqjiUyYvr5Q3t8wcZXsXy5BfBUrYn3b6O0YGoYZR2RMQ0qupHZo
HIvmT+j33o0uCQ8SonrRTeDizFGBSWBHqjzWNLFck9QONeRagtQWLmMttSZm29oE
ZI4lYJAKIvTS9yhvXdX+hFrr607ozcpgv2ciKg3MmYvPOfiFxdQ68P8QtjVtFkSy
Hp2b9KuiEeAHtREijjT0Fz6HcxuwVN7R9y4lvBbJWk9bMvR9euaJi4+cLjGAKEcJ
u8HVCjRLsYLxY54R1wPjrLjE4wiAwvNdpH1Y+TYW0+IhEffe9Ot6jW5FYho/SVKZ
0J6GXb5GfMppdU77371bsK95ciNgLk11j4I+5cqVMl4qbrK8MNTJbh7d/+Y0rdck
52BIjLiDl32uFyR6x26smtidujyjacSUT/6/0kma3zwxzA4Vwc2JoDJbFEjk9gCz
VvpUbSXhO+xYMaDVJe/JXr53TrxxWdkT1NJnafkdvtJRdUxH7UTMO81ByQzo63TY
K/crlylLt0HznZfP8jbTjoeif4wXJ7ySj7tT+8kMxBNPaPZy9TIFA0Be1PMxJ32m
Zc8sJCtci9QwHKlRD7PYbLoUDNBSBCZm8tTSmElwxPXOU/2qtylXfWh7N6JxPEhu
X2AEj0cBko0721coN6m4+iHiSfYVs1lwMP07DXAnpzLFhXL0mkLxRG+fpc/Sn9Lt
zBRIFY6P/eByby0T1mEUunWU+2qS79gYsCRIMaZAw9RysUeDpDjTVVxN1+QXKZLU
QFllau+9PhkSkKABNQhxQjKm3hFOaxt5p24XkZrTg+zb0Ie+e+Rxc1CmKB2+pWFa
8ljlyeeGBgNKoTS/Xk0KVGRPiFBHt96GX5NTLc9Xa55AKxNJrWdh3JwfxjD/b4F0
NM4YW+sbfn/mzxU1weBG70+IgKj0h+bKez+VcYayLxiHuWwgu/9BNX6EdBssTsJc
pQvzdAjjK2sJyskLDbL55CUswYYutie9+/UCgxwF1pWY0FDxFW6PWmnOKh+cVDG0
Sj9ZGR2joIi/OOjhiJTZNYxG+pe9OquUNOeHf5ku2NUjOzYbys8F8OHDE+sNK2x/
jGSOIoMrUUv6250hqV+2k5fi9btnY+DD6D8+U8okO1uOtSJBFQTu08UA+3+Um+t1
2MT5TjdLNDuOKc6Vi6kdT7dV5PgSc/qZe9A3D2CIgT6VFqIGy2Jenvd/nP9Kr1t+
pHHnoarG+ZUj0iutvdxS+/wDfwy2l0h+aggHwgS7iFlq05UwzLTBoN9M7+WXD9sA
PouJYIygkIdiwNddfiMnNpdsUq3+TBOSS4nvpddNW6dhjDsjDrd4bie6FeDSvohm
PAP8f+/gpiiN0mZ34xPifRG3IaKMi2uBYiHE9D0WpzjuJ84+Z9Rf0KQRN4LGoTG8
oG3x8NasvrzYZRvgUcIxfdobV+83W+isHCavAblpdKQkoPwm1ZrHtEepUteZErWl
o99DcjH/pHCRGQJXzn161Uk84llAMkonW1iywXQHXUzCkeNKvweablp+qwtd3N8S
QXxp+XZEWXcLiDJrmy2woCF9xUPxjB8xHjayGLUpRtgnyYsW8VHdHMwngzydjrEJ
UOGOvLg5PS4B3DvcFjML6vw42FbgZdUZ8iVaRuu0JYUh+f3aoMQIT+BMcsLEJ5Yo
73sF9EqHxLALSAjYfOI3t/hE00KPBE/BPXLu8HMQxOWbWspe2Xriqic5/UoRWHkg
jEZioesY12sd9Ex6Q/Bgtqvby9au5u2cgp1ZQjP07RVVCLavGtkB0lSxJrjdEW7D
0rgesKEn81Wc52GW4ZlBFzeCoFLuniyuApTsDh0SdVWfPHpGhWRvEaBzPJ+40IKD
yrqH5hqp/zXs8f9BcSC2OMELASIOgTjQAdQxmFCOodFoZBjL82RfYla/FalSmy1m
RZohIplmYYtex+aLCAJ6DHi9vdHudCt57NduzCk3MQgnB5mt3m9W4qAm2yQetKUd
OZEY2OpE4T2AKphRZL9ZiJrstlhhbgUyh8DUaOci9/fX3AmxA38jOBUeHEVryP8B
pcImgNxEmnRT/YiETeyFsZrTfgBStRRfdOkBTp7tJHtY1Yfzqh/JTvBkIQW8Vavu
FtVI8rUJRiDX5n+7dMtrrF/q2IEV3OiyjO7pc7RNtmVH9XhRfvjZIjsj12Ru2+7U
Jutts8pciyRnMxPfx8lxlrAvng43UpXRHEd1cAfBhjWCbve+6iQjL7hsLx6ZEKTX
yh//twrwR9ADxAJptUx9rC2dHIzTZXBb1DiAXvcquy+5rJizxsrS1j5JKusaN9e1
+U1u10LwAom8CoXzxMgET3kfHw44Rw/ytbAWHGFfpxRjm7syrYne5a/oPeoTIqU7
YWdlOFJHNkF1QYZGg7VBo7YLFAZH58Fl286e5iWS/6+wZJWt+/u5ShoPyjh8qp++
hhojP1FrymFXmCdyMVI7/6x9lCGx/jFxLbjIgErwLnnQoVGBqUM6Lu49T6rTTGFO
L8zc0nVKYCtFn5dXW8aaekqBdK87xlVpXQ6vrDuAlGtuyveEoQqLPFePsDW3+XKY
6uRbMROezDxbklHCourMCvQQJQocW8vOfUEZiKr/fv4MzmKZEU3gm2V3YhT4DrpR
JpmopMUSQfehcKY9jHjdxJrYQztuM7csoTKPBgexSxvdYYVq9q+xA3dqpULEW0UO
MXeITb0XUkiaZQUQoBNn5FNx+qbKEZd3luWuajh40GKVmWvP2aUSUrWLw/on0WcR
Ia9Jz8bpxo2KpGKtUTSRkXgdapz4QhlT8NHzVYN25I6O2XNkbbHuu7e04Zt2fUAJ
RBRjj0ErS9ZurzYSwtBoJqV9DIGhn/DkLv1fNTbwkqxU1uozCNsnMrriNZxiI+h0
mrBuzt1v79kHyQdh3IMiPk0+MdNymKxqcs7JzhWLu2kfbEMDsP0CufRGemiEZFiM
IW7fkuAdeoZTCWYhWuuI06HU3PsMauefg7cklE/e/z+/q1+6+nGKIv7nwEPdvfhE
4TX760fWa62DsVfISuos/dRSpfVUqXdx/8ZdQzC+mK2wCsQmUz50h/xr2nK4pAsK
Va8fxYHDwp6VSJDppr84eoJIGiC8n5mziQPnooyrpTdSqkb+Lu2a7y7cabIgwolJ
CEt0bZw+1tf2sFLjDqX0uDnqdHXmAgr4KreThvoMcveS4CgUEkd8UrTVim59X05h
vR8IxofpeftnQz7nDryFUU3FSOoT0ks/kZsA5uPtynAh+RsJkUoU2DXyLnhr4pzx
5Rj5VWgKoBXv1QbNzR7T168Lk2AE1AVxsE1FaBlbZzax30MU+XAQTlPViysVSNdf
3FIcO56AlXm+x1C9rI1AWzl1s6RPcsTQ0ULiCbShbjtw4+QELhmDQwkLqe5EFgR5
U1l9ZqKAmMfmLEQmwsz+d60NUIJd2lPUAbiqLeLy9KTWveJwCp3Gl9sHCErEhq+5
XkYueRgBsZrqhSzQyp7Za9Eaxsb1ZvlJ0bErfo8eOijWVpIwf+3mdRI/JBYZaxqC
W0jLT2xVekOFNA+gUkgTArz0Ba1XXB0FfrzuTST43Ai4YlvVqaYdWUxdXi+hx157
LTIYp2EmRqfCrZ0T/4bCDYEeRYrAQSA2NhLvSa3qVEj29znXUHIt+BpX1n1WmNHP
eYzY/BZ6dqXiot8F06n5uP3pWXi9O0+fEXMyf3dfgY6XzfQXyV4hjGssFPmG8y3V
8zEnnn9JtNtgxH82Ab75P9jB61SwnD9tCVUKZBHZQgI8nzrA6JuhGaL6LlVHLFyf
7Z1iMfzjvD/NkDbYTSqNLW0NNGuUloho8SoNDZjp8/1+CJRfeXsDXpxneIfbgw9f
40dLDEpG0C/bAVBrQKSeat9QYh6Wb2N2p1EoEcTcl0dVF0FfWob9Pux/SAzi7pI1
AAjNIRUHq/0aeL6ba8bmVux6tdfslhdw/KAqfC/xICzw34QVnF+fuy0LSAfjTrxj
2k441ngObzysef7ZPZhJIW/DFGBf77xooVpaEcx2y+QXOIHrv5VA7v3XjEV6cTIS
kTqX1OK1OaC64MtGuJzAQz++NOHlXOYh9qCTxi1hgejh1yOTWb09UyOiKxJ5Dl0w
dyNJvuvEZaJ3HVZDxX9eZQERTA0VXLrG1sKMCQNakc7jDII2svzjrz9iktrUmI/S
0+UACcFogrrJKRAyQ39mY6InphPA+PzMIVS2y0gd9zidTdXpdT5ff0W4GOfjtued
kY0ySj/bWjzKRu7FZmCnsOr0lBFCbj62j59ag2vEtIE131O7QzmVrGSrI0iGdwlB
aQVVYqfHQ3YJAf8SjG43nLkewMM5hjSvBm6wL9FhXYZzwec6K+suFgAkSgc72QsJ
YxuPWnP5Sdmq8aboRkCDwmz9ERgmiEhcPClEhdsmHKuIezknAZ2J4uyELU1AQmdm
NSqKofvEPkIaT5a5cn9M1Ak28DflJh6GDRHSz16GZ6egmR5P0IKGEWPNjTGEYQ0g
+yVKnCg6lp+wSNXf3/jQICUOrASDk71C8v5PnD0GbB/QcgGUFsFuK5pTIrf8yIMN
sce1dQhF/977MnfxNKFHgsxWHKKs5bQyPZkeKWNZp+1oU/+hnXuYOXLkN99NFmnJ
n6QO+N9J8wQR8wYBIuvbRw8/erLmZ0rGHEJcBAXUAi6TTES0I9uOAqUVW/vkq5MS
ssPLsw30WBnSCUf5caIbCPa0IIpAWxG6AT+yw8Or9VQcxk0HonrJh+0qE8X0jvHH
ErfczeklBx1SuDDqgPZu3ja7o/N4cQwriY6UdeyCknXw/qX5CROE0zTE4tG6xTKp
uCOCklk/YndVD5rThXljYygtBLQdob6XzNh8YYA6fjPIpIbE0JZyUeqYTshqDi5q
2DWLU2AHppqxqSreV9efHKljkEp+bdjMzis/PPWonVR0UsGkji/rXduc9D+ZIUCb
NB2WPUykYi8T5QawE1bB52T2R+U4qBE9X2FFsZ7uHONkj3ALKamwysc0kszWBfUu
+Bd6AieD2mErl5Wc73NH8U6dgRSc2rDogq7MsPHrDRsqYrYXv3U9zVX/Lu0YK3hH
xEooci433+CupdvhsIp7fBPimDlg/V5naeZSZbkJ+DXEnObVS5s513Szj4f4Wz/f
kV8GnjPfePpLJwJ0RdDvzXsKuJJ2WOXbnX3pwbJvm/70KivrUcU5Zuk4Hwk69R84
AOQWTx3SQ/FMOaFxBYOeQWtguwkuWGNsgooLjvF1r4oajhKbDBacKlAbxQIRIva1
BpdzZU6IKa9oGtPa4RKnrNVs1FN6d+YwRzKxHEahrZ/812nBnRUsGEC6nARml/q3
UTEUIhtgzVjFdNh0Mksw7evTqgEsfpmJ7QuORuiSfm+Jj/LKeXS9BJSuR9Ke+b52
AQDCPR1Q3FrF6IDkwfo3tGVETvtvJZvNoAVDio0AugnoMysNTU7GbdxsKH7uZ1gE
/+nxBWqeA4d1riAVewvyDtm0JUssCUudFMZ4KTlRGrRgMSv89PEBZecw+RG3jRCe
oGmFqNHoxv1lQxBCWKfaGs+LcWSwuNUM7br/hwMpQTgl7Mkv12OYQiB44zaEel/o
c7zCPlDXgJyaDEutcNweRR0ISLrldW6hPI2PoXP36/U9N4IatQRq6V0fzgZ/k+QC
jmnIK98WenOZOGilShyEeAgTave53GcpZ803DfFpjxIUdUHvhVH6+hvpNHR9MNAO
kCpUy4+SxhVkCnr5C56DauA1mM5oefisfGJ+hdZSHqLv+0hOZI2anluSHug2pk1F
s6KrjvMtfkmik2YhPRzYvtun+id7gKeP04/5Rt0u8skhih3Mz05DdkvTtN2BL9NF
Qli/jo3zupeTAGOZ8vB5dwO2yhQlA65d0rRS+NzgpbD6facz4c8gz1qwU/Io9kDX
ourKZjua3r/ztQaJ0zyJDy+EOos3sW6DEdLk1MttoLuNnL6ovCR1Yzxq55ObtaVj
uRwyvyV6g0ZEZjZsEWXsvGghO0ZgCixkIrnPyTNkIJXzHgg1RCbTpnFm9nOUyOyC
h0dqDcjoz1p2a79AhR0RhLdjE45qjceoc7X7GA2ux+fKaXyuBipIpUDaQgs4GNSZ
4OAbMyJmZR+g+usPjiS4L/h85UicqAmU+2CEoRKNrM7xy8FlLnPLuplNTfzL2mcu
uBGpRXgJihWve1HA32zPi5Rn/TRWw3Wqc8hq6s8JRje3G4jsn5YIT1RHwd/CGzLH
0M7Dn5QvqanX9Bq9H14V981BMmB2J5DRmD90Egt8fGQ+iLSEn7gfqwBCeL/sXnaM
5erRLCa91J0VpybIFSX+gXTtUIb3Ow87CA70IxcamiEtFaNka3NzsRfVG1OwZvJj
t0/n0xHuhUjlpJ2ERdXQcRxz6BBvRvF+7dYjq2bbSkjWmmLlKfJCWN7hvFhpvYBR
XCcVKV9EOe7vUFDtcpN8bwjFTPXbXbVD7fziR3KdH96hH11Fb3W6fV2RqBKtGT1s
ruzpMsYnu+QDCqpSMGmv5MGZ0nyWenBBXsmeBQ2S7tB6PTUL0gWjFVCVfm/72mzo
HIa2RcMWBXZuqrc679d2665qakddlzBWLjKygEqe+pHj0pbu7qc4ZSv+4VRnKvtK
UVk+PgMgYaa0gXhAKNyzj0atlwyUCkqIoqdUed4wZlwXmfJrXbop8zmO3nrsmRmL
ng3rt7dotdwnfnd1NdU2mWi0s75EW/zdN8/CWparRA+bymBpuDApmXaB/pMytnOQ
zUZuuI+2bfcYQzRo/WPi1h0AfAZOH3/rRwdZSq+oQpK2O2JdmIob+Uh51eEpoA0I
9hpKGDhhl6pKXq+RL0r6Ux+IZ0loL6nZ/0wc5YP+Il3T3t6mGEJrcmu8QftIFBOU
5M/JOzXP7ZwqozEpXV55hBcoGr2vOIYv4scn1w9j4lv4OSMF1sW24PuCW+H77wHR
c1AfSANS1KxXl+mCZNX/20QZwWymCyZ6RYfYOoipy1GrSwZgdbx5yNzMg6gqbDAG
gqOiZyGGv0FZTvx2l4KHv1wTtJ1oUhgTkm/WXuKN7h6bk48sVlU6yDpDqeeCzeej
iIyw85jlz/0452UwX6iweoL2yHlfGwcgpol9wvj/u4ZW9MPvxb9C87Y56KZba/m+
FCM8gTjjbsZ3QdLmodDvvwrfDTK9T9iaCBFRa0GpSrSHC0+qW0/8V7vVXR26sJpq
DtvMAi+1a3AltLOTfD6q5sKRP7gfc6tnaKIePnysGromkH5DjZg5ez7gR2R18a6c
g3OtOGKD5BiwdPjBpQggLXwP080R0Oafidin4novXRK0H04vGM0rGiAoyzvRfybS
w9zeYgphWFVhd7FuvLX6bXr+85djA1vSn06OE2F77wrx+2Vvxx/v38rzCNbkTBFD
qzzoAeMyWzwRM4jBa/YVGh5gOtpkezZYzfdXsp6aY90NCP+M+JztQdrFtaRjcTxP
g/b9tuNfsnnszhy0wHUrOZ0aWlxtC3QykgTQHj7GBY0fUO2c9WnMSi532Uh6aqLs
pQwnsoH1VOvZ2JfrtjsPZmEIBrrUYKvYZT53nnk6Hmp0vUVB0mlGhDX/H/LMB6KK
Hvihg4rso0lBFraUmK3yPb572ToCV7QeWZhDn+w7NA79MMAHlN1zDceaUW2SQII7
VJO7b0ay/l7OVKIVYnC1zZkHR0rgvioLPyT0ldUHkPWakuUdVRNLXfCselvQI7jf
PlMyxK2uj+q67a1MjYOkxNHhsLBrKVC5fZXn7XlEtn1bpg1BK6y6OCGiDP1hjY6d
iY99xfxreTfsUabv3oIqGWa5N3bFenGEDFD2oOvgm1cA3HidXky/z7qhkWG1xs/p
3MDSZekli6ese6yURflCcQ5Z2G29G93zlTamoXfcCkYyOfpPXGRQHdWt3YzuvkEa
tlaT9dlkGJr++ts+RZD5BPgsEK01krI7Ap+nBFD8ty1MOqOocI/3frL60mocwKZd
20q068EAaqcxsf118iIUldAfdCAJl/xNWryL4+Os3tKIz0iHBus+1coJiow7KLjW
sc/BVo9iuUxRIIKLbUwPm7BJoG/U+r4lmG/bS4nCpJlWtmMpvfepE2C2vrZ/ebTH
iQGJ2p2S0ltIDCvHkkdDgJY1DjStbqft6Cco6ekPhkJGe5fQhKZ0QjocEBY9umQg
Np7X7fq4vlp/0Y34fJo+kJCkDWvlYG5lPrKTxeIYiRuw+kvPz6Z9w30SJaKHjEoa
OPNZCPngaK7+H6HGf1SaICJci2aDeUM93r/FE/LEEHfrKVnzrzRalv0HbNG8XNVc
OvSP6WrxaSzp0a8SzmAMRukgxSq6SEruLYmcE/4lQJkAhmqMr+3I84LRPn9t79F2
tyyHY8F20L7QFpP4qTLLt6w6Xv+67ZtzWb9Z2hV090QF8fMhRtAbppBAal8XglTL
JM8eMTUNVRItHtooT6Q6sap/Wnzz4gd5/l7cfCtNSDgqPqOGs3vODPg7k587g72p
TRClTNhHLVn9XJ2H6UZzgz4XlbM2E0PCUJNJGzQOuJVv/0ztFcXrnIWyNBoYyw5s
Eg64A4FyDvEYEV5tqXWWeF0rE7cHMIKcl01jwM2dw34wCCNnOZ124IYbM2Q6yNG8
tPUu7DUEWLVA86jLYgZeTTX6PmPNcdIivA2xm2OqOfmAVmEo0JiICywqeu9S7xI+
mWVJtZ0YpvA9WENXeSRHL8XM4D6tRHbnbSRvKgE7g/o6lWvMN8k4D0bV7MOvDYT5
yQOSKDcpqwrbgzf85fGaB+iI2igzikfsdst/k8cCnYFu60zHk+oD+MuDp5g3hH3R
OPeyohOR/XmQ58JHixWIHwlt4TCkRrDRdrTVnXOUakBwcU2vFWZp1GI006En8+b3
ou05LdZrzas9dUIvLw6VH9rWJj3yhxOzIQa0xLYJMLOFYiwwm9GU9ewWcWTuvquF
C/FwFaHK85w05a1qHKdYk3bri4Rzx8qt1br3iwqi3hKj8Cajwy1p4lXPoCgYRCC8
z0CiXi/YaIS/TzmMScvLrv9stYthJvlBeaRp59Yru03MgmiSkp+E+OPZMirQ/M+B
iYVxVWwjLrzFzIM+U4BoV6VPO1SjxH3SK8whK80fsoY/N4xZ4dw5UyNtV58qtAnP
LmrvEIoRm3I6WTAnawomXB5qIjezAyK/CEkTA280bIWceiKHLRWFlvR8/2qkdrVW
K4+ko8q5YWNgbrqpf/3wVNTI5oxcxc2ELm4J3BUZLIriuKBopi8T15BCrurpV4Me
VDb/8e0qVuNs/DXWIVpqQ06jOdvuwczdJSjG+X5H4Z9ADsTnzBvDY0pJxKvBUbEV
rWPah6ckxPVySFCVyQPJ5gmI2/cbTwp/lbHRpUDmpoiW5KlxVHa8R14zjIctgZ5d
OXpb7T5x30aRdpSnyM4s4AS79wfwpDz/sWhJQm82rNowxgbh+vEkPVp/7DXeBZcY
PixZ1Ae7fAEz1RYsCdkcCzXsw1xLssuoFc2Pr49G50P2O17AM8DAB4ku+5LJy1SF
Dq8h7vxMoqzSI1gpxwdnxUqCEJttf5onJfR1udlyJjzJ7x3xgIbxP7x6cFPp8NaW
QShd6czaOuYv86Ci2rX9t5E90tW8IFT4+cLsK9iZxwEzovqqL/vZz6TwHywtfOjk
U7ATqznzyU4IZ6jTxsW+l7uz8P8rDO1O2h7a6Okmgn9TevktQYtVZFF6QWaZg1tq
3bZ/WBYg7esyKeOU9w0531ZeIxULIkJi6QZd4gbnlYUsNKOlJljLXCzat7epwrM2
evVjQ5stgFDDeqLL6rCeihReYZYAC/8YZx4zBs2TeP1F1IKDUU5jeZmulHUUC+TB
NxiFFbE2OZX4newqSZF0Uw4HvtHln12ut7xTdQ6Mzby4SIFQC2dBZpc+IIgtQCCK
deb6eoWJeBbfXyzxsolyPkb9l8L0JuLhevEaLoDAduBpczRUzWthBQ+ILe+JDJL+
z+YNumwzTlPnLVk2nFiyHcrAwaFSDbOYb2CdxmqUChUrxVTJW9f16W8K9h9221Ov
IouuNvq6NC7f1bT81vLYUvHW7bo3Bo5NPkOtI75MvISHaTSSh2CPb5xZOAi3R5S/
QttdpxTj6g/HcaYzFzoY0c8Cc0CAy+Qc9DKHBhxfHtPXxIYSfzY8MDkIGcNWmaDR
ELe8A6DU5iVZ3RTGFonk2HKYkLl9scI4vzLrjf6kGozh71wIjoyqJZZNPFBzsimO
iCEPBy/PvPxlCGEU1TgJsWw0kIttHucq2cYxTwQsNF1OSDu8PBdY5ituRyKVRlxa
Myd22rck2D0yJaCSN8w5cb0bxo0gfHP/GWezXNmOLyu/XwkvfE8yCTM21L+KsKfc
9AqDwuNNx9r2wlg4ayL33DCWKMh74pFnrbz4KbgNN+HS9irw2kbsMtSdKmQGzdo8
rx0dIkIW1WJZXvSl8Tux3i3QfsjKVUV6zEvpSBYdGRhpUNFND/xWYFesrCNhr83i
sYK/DfmDG0lARrJcc/rZcDHZDnInoily2lu9TenDKi6pVdV7uV3yCY/4AwzABG9H
USgdnXDp1Itx6/xvrUY69X/lIVzNgrViUZTHw7/Wlbay6HmpNWtdDgquF0ssJ405
oHFyrAuvFzzzi43B7W08LerHrH05T+a5b44gJk4xNPLOhwE0UeOX5nqsjFP2FQpy
T1ehda1T/GdSIARR+NAbyVt4MttzcRkdmn9qPse3O7d8Iu9O/BNTs9Hxa04ocS5Q
gRwN3t3kRH/kupyf0xQfzhQWOO2zyaAa49P9w4xe5BzrLTAzR4a0xDqQ+71cQmV5
oxLxog1U9okRUXsoYWM/IZFjy+ssAWBngEJCH71IdUSbMQM4vjoQBFPBwraAYBpx
2HPq7ib417W6mrGqJw+m1Dddo6cY6EniIWxa1Uuetjn/Xda0c8ic70n57ObfTdQZ
hS8VKjaJUQMdpND8FJowvGI5cH9rX0/AQFjd2/omkO5fqNkWJIYoaqYCbzpI0EYj
KymdqLniLEFlRatQWcQs98QdpyT4N1UqWm5U/k+TMEVy8YQtPsp6LIHd2iBQavuF
f9xR1/1oIDManX0ZH7SdKobBv4gvJmARrjaaJFzSVoXn1beRxc03yumRAyl0Q5SM
RnZnGPwaXgszEnKIue9wuvuopQ+C//fWvFazizUJXKSTZaIhx6V+nselAj7ahddf
SZa/WkDvzsrbuSV1yHQIUCRw/ZPSM/mag9oRfOEjz/hddlY/VgpNyteGRzaEKNFQ
bZ6PobfdT/KXmE0dcCwD9wQnZ0AaT/foBnudaP0jV/q8olG55tw24pm1VeHR1fIM
7aeMXCcY4vAlIllUEanoRV/K2gUsS29w+f4HeZgTWz3TLy7nefTGZY9fcaRLVGMe
bhQcrUhY1kmakVnFjnNda8YBUw26NoESereFcK1Gjls50eHw2uzan/LuimWAyuXw
kqBPriiCpdo/SZMQCv/DqNiIA5RrrewX0Woo9EafwPl9P0036Yo+5WQpPcVNRaOe
lZ2bembjPi4j6NjGZmTCuG7hHTMOOzA1pUsGZkSymDhxLVug8qOT5SJ5jflKOSqe
Ar5Xnd5rXS4wtbQnoshXtEQweeSNkgrd/hx2erFbQHXfDOuFNfBkCXor3Pmm5r88
vlqyzzXX8stxSM4VDNs2bM/3JYzDprhBEK/04UWxBu4ktZl+t046emRZ9C0FDKXW
NIsOZfLVQhI0TgAP7v7xvY7+pTxW+SrAr2xeF1jK08j9iBNjFX/06rx4ut4VVL7F
x5ms0mIqdLlAfSiO54BULzqGoqkkwk0ZeRuYWOVeTn0xfRwxVF8Nzz5kpwy1xIDS
Df237Y+NKdR2lhn7Jy5EW6zyVVe5fFhNzneVfmeEEm68ZgsGefT03hR+3Z+hcZne
y0Qutb5VfCU6a9jdNLny2Us+gYaStKQ7GG8ByIHOnQnik3EFOu9o0KUHkD+wzLXp
qd6B7FZQc1n43qxLnUFIFRs8JepVdB/O7aUehE0mmEHnhlV2/F7KkLKuGQbhpBO4
k8Askpd510nQMUKU4t0nLMXFNzPQj6FSTJ9f+VXOJAHczpUysDXDf2owg9Ya6TMN
2VvqsKZxjqAOI32+G7cyQWFqaTI0dfyYc90X1FoK1w3IIbB9x/xh9iguWdBOuCRg
eIyYeQWK/BHgH0X1NLOpTU/YEi7f5KKQXmKhvJ7YobYjGlsGtapnX7D59byeE2Fk
eQ5Dw0G2R16M0lMmRAzIuRL04BwT2Zj4+GPc/d18Llaq8SpV5ko5pwhjRvFtQ70d
EEvPanKw/dqiQtiIih08TWuJyh33U2hB+xn1dyMUnOuS/Zt+SNgJ3hwpvmYP0K8n
z2yhLsCJUyXHlk3HGr7ZskuePQmduOAJwUufT1sLsPjI85tI+UK9yOPyw+3cCP8P
aURAZtIfW/RldtxUUr9GgySREuaxYz/T0yMEn1wh+8v5IyZE5MBMfjbJXFyt8gV2
slxRwlmjKWVvu2r3LPqtUy8kN/4tabP86nKCKJHm7NBSeM3ww8WQjy4VKz3P41d7
ajw1jEQvH9TdTYZkaiNErk7uLfGcNzKHnbz9TWbxpDCczd+d+vq+NfBOQhHqPKJ6
frYQfXloWD6wCa+2X53bV1xWnuYMDHxTWdMdP8pzHB2i6cqH/ZPRtjpG8nvD9N/R
ozgrButo9tbVk9497koIQo1LC0u1h6aFCcjBMONWx8N/o/Hm9vLpigO5TpPRK9do
5z5TxlBX4JWQ/rX8O9dtmqCllceucxLY12Fs2O/ZUW8nnndF4KqvPHV+Aweo59/2
4iY9fGbnZbiDz1cuutCe65Pcz9Gct3YmA1aO78Q2NAbI6Z2wiZ491mUXW8lvYlQF
SGmglRH2uIXg21gRMKqA70V4JI8gxjANXfaJhsYIavOp2oxLHrN0Q59UaIemhwOz
EUC94AyN0eO8aq3uEyR/ElI2eMv06WRTTvvah9xhB5Nj8CoLN+5QO3DTAXMxymfI
T0gqgBwSlgjPYpcyJ+vWoEIWxINPwjjMyMjDlAq7O6jCOCgMnwQs2uypiTzi9wa2
srIKG/OKmMVA7W4fYj/k4iOjm17uejT45jtDW27iGiohl+Out9k0mFtg5vYa4p5o
WoZKUM0V9WBfBMbDU5xS5qjKiGTiloTYzjK69uHR7EzNY3obxxruAavducvmwtsG
E+fq8hmsbYUOtAz51svzm0+BTdyCo6IBp+IfeqrTLbuKKzMAwtJjOL9BD0w1RsY0
RExJGkgUZ+KOrxPdf62ZqZGEIvbFhY6KD2zpDfbpH5WDFQYrzFpDk3OPQom1MdyI
dDgkItZ7FQ5WPaMpxQCztl5kM+fhjujpqomrzuyBO4gxZ2UAeDWP+J4IELVRN1vn
NEKqqK2EASjySzsfxOpTb73bs1vUO2R0FxzfPpdDssI=
//pragma protect end_data_block
//pragma protect digest_block
qPkTH/xalnqH31JZh7Qb4IhJ4Dc=
//pragma protect end_digest_block
//pragma protect end_protected



